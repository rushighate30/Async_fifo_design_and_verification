
package trans_pkg;

// `include "enviroment.sv"
`include "transaction.sv"
`include "generator.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"

endpackage : trans_pkg

